--============================================================================--
-- Design units : TestGenerator(Timing) (architecture)
--
-- File name    : testgenerator_timing.vhd
--
-- Purpose      :
--
-- Note         :
--
-- Limitations  :
--
-- Errors       : None known
--
-- Library      : BitMod_TB_Lib
--
-- Dependencies : IEEE.Std_Logic_1164,
--                ESA.Simulation,
--                BitMod_TB_Lib.TestDefinition.
--
-- Author       : Sandi Habinc
--                ESTEC Microelectronics and Technology Section (WSM)
--                P. O. Box 299
--                2200 AG Noordwijk
--                The Netherlands
--
-- Copyright    : European Space Agency (ESA) 1995. No part may be reproduced
--                in any form without the prior written permission of ESA.
--
-- Simulator    : Synopsys v. 3.2b, on Sun SPARCstation 10, SunOS 4.1.3
--------------------------------------------------------------------------------
-- Revision list
-- Version Author Date       Changes
--
-- 0.1     SH      1 July 95 New model
--------------------------------------------------------------------------------
 
--------------------------------------------------------------------------------
-- Naming convention: Active low signals are indicated by _N.
-- All external signals have been named as in the data sheet.
--------------------------------------------------------------------------------

--=============================== Architecture ===============================--
architecture Timing of TestGenerator is
begin --========================== Architecture ==============================--
   -- This test suite will test all timing constraint checkers 
   -- (both with and without timing violations).
   --
   -- The test suite can be executed for different simulation conditions using 
   -- the SimCondition generic in the entity.
   --
   -- A listing of simulator outputs (assertion messages) is provided in the
   -- reference files: worstcase.ref, typcase.ref and bestcase.ref.
   --
   -- No verification of the signal output is performed since the main purpose
   -- of the test suite is to verify the behaviour of the timing constraint
   -- checkers.
   --
   -- The timing figures have been taken from the data sheet for the
   -- Bit Modulater dated January 1995. The timing figures
   -- are based on 25 pF load on the outputs. The timing parameter
   -- names are compliant with Vital Level 0.
end Timing; --=================== End of architecture ========================--
